module vgdextension

pub type EditorExportPlatformIOS = voidptr

