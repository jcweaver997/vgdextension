module vgdextension

pub type LightmapperRD = voidptr

