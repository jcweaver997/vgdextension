module vgdextension

@[noinit]
pub struct AudioEffectLowPassFilter {
    AudioEffectFilter
}

