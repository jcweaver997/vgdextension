module vgdextension

pub enum InlineAlignment as i64 {
    inline_alignment_top_to = 0
    inline_alignment_center_to = 1
    inline_alignment_baseline_to = 3
    inline_alignment_bottom_to = 2
    inline_alignment_to_center = 4
    inline_alignment_to_baseline = 8
    inline_alignment_to_bottom = 12
    inline_alignment_center = 5
    inline_alignment_bottom = 14
}
