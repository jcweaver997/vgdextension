module vgdextension

pub struct EditorSceneFormatImporterBlend {
    EditorSceneFormatImporter
}

