module vgdextension

pub struct CSGCombiner3D {
    CSGShape3D
}

