module vgdextension

pub type EditorSceneFormatImporterGLTF = voidptr

