module vgdextension

pub type IntervalTweener = voidptr

