module vgdextension

@[noinit]
pub struct AnimationNodeOutput {
    AnimationNode
}

