module vgdextension

pub type Tweener = voidptr

