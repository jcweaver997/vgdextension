module vgdextension

pub type VisualShaderNodeVaryingSetter = voidptr

