module vgdextension

@[noinit]
pub struct PlaceholderCubemap {
    PlaceholderTextureLayered
}

