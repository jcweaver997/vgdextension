module vgdextension

@[noinit]
pub struct ResourceImporterOBJ {
    ResourceImporter
}

