module vgdextension

pub type AudioStreamMicrophone = voidptr

