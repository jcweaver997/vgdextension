module vgdextension

pub type VisualShaderNodeLinearSceneDepth = voidptr

