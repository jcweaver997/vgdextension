module vgdextension

@[noinit]
pub struct AnimationNodeSub2 {
    AnimationNodeSync
}

