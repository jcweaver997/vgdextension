module vgdextension

@[noinit]
pub struct VisualShaderNodeTextureSDF {
    VisualShaderNode
}

