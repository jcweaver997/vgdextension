module vgdextension

@[noinit]
pub struct ResourceImporterScene {
    ResourceImporter
}

