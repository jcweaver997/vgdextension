module vgdextension

@[noinit]
pub struct EditorSceneFormatImporterGLTF {
    EditorSceneFormatImporter
}

