module vgdextension

@[noinit]
pub struct HScrollBar {
    ScrollBar
}

