module vgdextension

@[noinit]
pub struct HSlider {
    Slider
}

