module vgdextension

pub type AnimationNodeTimeSeek = voidptr

