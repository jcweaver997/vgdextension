module vgdextension

@[noinit]
pub struct Separator {
    Control
}

