module vgdextension

@[noinit]
pub struct AudioStreamPlaybackOggVorbis {
    AudioStreamPlaybackResampled
}

