module vgdextension

pub type ORMMaterial3D = voidptr

