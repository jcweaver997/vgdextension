module vgdextension

pub type EditorExportPlatformMacOS = voidptr

