module vgdextension

@[noinit]
pub struct TextServerAdvanced {
    TextServerExtension
}

