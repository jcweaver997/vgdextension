module vgdextension

@[noinit]
pub struct EditorExportPlatformLinuxBSD {
    EditorExportPlatformPC
}

