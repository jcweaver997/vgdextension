module vgdextension

pub struct LightmapProbe {
    Node3D
}

