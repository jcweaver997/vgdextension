module vgdextension

pub struct EditorExportPlatformLinuxBSD {
    EditorExportPlatformPC
}

