module vgdextension

@[noinit]
pub struct VisualShaderNodeParticleOutput {
    VisualShaderNodeOutput
}

