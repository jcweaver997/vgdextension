module vgdextension

pub type GLTFDocumentExtensionPhysics = voidptr

