module vgdextension

pub struct VisualShaderNodeIf {
    VisualShaderNode
}

