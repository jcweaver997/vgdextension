module vgdextension

pub type CSGCombiner3D = voidptr

