module vgdextension

pub type QuadMesh = voidptr

