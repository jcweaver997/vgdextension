module vgdextension

pub enum GDError {
    ok = 0
    failed = 1
    err_unavailable = 2
    err_unconfigured = 3
    err_unauthorized = 4
    err_parameter_range_error = 5
    err_out_of_memory = 6
    err_file_not_found = 7
    err_file_bad_drive = 8
    err_file_bad_path = 9
    err_file_no_permission = 10
    err_file_already_in_use = 11
    err_file_cant_open = 12
    err_file_cant_write = 13
    err_file_cant_read = 14
    err_file_unrecognized = 15
    err_file_corrupt = 16
    err_file_missing_dependencies = 17
    err_file_eof = 18
    err_cant_open = 19
    err_cant_create = 20
    err_query_failed = 21
    err_already_in_use = 22
    err_locked = 23
    err_timeout = 24
    err_cant_connect = 25
    err_cant_resolve = 26
    err_connection_error = 27
    err_cant_acquire_resource = 28
    err_cant_fork = 29
    err_invalid_data = 30
    err_invalid_parameter = 31
    err_already_exists = 32
    err_does_not_exist = 33
    err_database_cant_read = 34
    err_database_cant_write = 35
    err_compilation_failed = 36
    err_method_not_found = 37
    err_link_failed = 38
    err_script_failed = 39
    err_cyclic_link = 40
    err_invalid_declaration = 41
    err_duplicate_symbol = 42
    err_parse_error = 43
    err_busy = 44
    err_skip = 45
    err_help = 46
    err_bug = 47
    err_printer_on_fire = 48
}
