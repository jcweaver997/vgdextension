module vgdextension

pub type SpotLight3D = voidptr

