module vgdextension

@[noinit]
pub struct AnimationNodeBlend3 {
    AnimationNodeSync
}

