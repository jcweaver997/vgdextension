module vgdextension

@[noinit]
pub struct GDScript {
    Script
}

