module vgdextension

pub type VisualShaderNodeScreenUVToSDF = voidptr

