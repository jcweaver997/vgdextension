module vgdextension

@[noinit]
pub struct SpotLight3D {
    Light3D
}

