module vgdextension

pub type HBoxContainer = voidptr

