module vgdextension

pub struct VFlowContainer {
    FlowContainer
}

