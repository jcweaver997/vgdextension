module vgdextension

pub type ScriptLanguage = voidptr

