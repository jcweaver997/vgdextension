module vgdextension

pub struct Tweener {
    RefCounted
}

