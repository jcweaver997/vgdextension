module vgdextension

@[noinit]
pub struct EditorExportPlatform {
    RefCounted
}

