module vgdextension

pub type VisualShaderNodeVectorRefract = voidptr

