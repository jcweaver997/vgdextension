module vgdextension

pub struct AudioEffectNotchFilter {
    AudioEffectFilter
}

