module vgdextension

pub type JavaClass = voidptr

