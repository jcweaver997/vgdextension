module vgdextension

pub struct VisualShaderNodeCubemapParameter {
    VisualShaderNodeTextureParameter
}

