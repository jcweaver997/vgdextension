module vgdextension

pub struct AudioEffectBandPassFilter {
    AudioEffectFilter
}

