module vgdextension

pub type AudioEffectNotchFilter = voidptr

