module vgdextension

@[noinit]
pub struct VisualShaderNodeTexture3DParameter {
    VisualShaderNodeTextureParameter
}

