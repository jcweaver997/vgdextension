module vgdextension

@[noinit]
pub struct VisualShaderNodeVectorDecompose {
    VisualShaderNodeVectorBase
}

