module vgdextension

pub struct GodotPhysicsServer2D {
    PhysicsServer2D
}

