module vgdextension

@[noinit]
pub struct VisualShaderNodeSDFToScreenUV {
    VisualShaderNode
}

