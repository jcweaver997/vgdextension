module vgdextension

pub type OfflineMultiplayerPeer = voidptr

