module vgdextension

pub struct VisualShaderNodeRandomRange {
    VisualShaderNode
}

