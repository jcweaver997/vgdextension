module vgdextension

@[noinit]
pub struct VisualShaderNodeTextureSDFNormal {
    VisualShaderNode
}

