module vgdextension

@[noinit]
pub struct VisualShaderNodeProximityFade {
    VisualShaderNode
}

