module vgdextension

pub struct EditorExportPlatformPC {
    EditorExportPlatform
}

