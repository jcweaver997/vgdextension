module vgdextension

pub enum ClockDirection {
    clockwise = 0
    counterclockwise = 1
}
