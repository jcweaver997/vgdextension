module vgdextension

pub struct MovieWriterPNGWAV {
    MovieWriter
}

