module vgdextension

pub struct CompressedCubemapArray {
    CompressedTextureLayered
}

