module vgdextension

pub type VisualShaderNodeGlobalExpression = voidptr

