module vgdextension

pub type CompressedTexture2DArray = voidptr

