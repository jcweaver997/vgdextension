module vgdextension

@[noinit]
pub struct VScrollBar {
    ScrollBar
}

