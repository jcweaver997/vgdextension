module vgdextension

pub type EditorExportPlatformWeb = voidptr

