module vgdextension

@[noinit]
pub struct ResourceImporterShaderFile {
    ResourceImporter
}

