module vgdextension

pub struct VisualShaderNodeTextureSDFNormal {
    VisualShaderNode
}

