module vgdextension

@[noinit]
pub struct ResourceImporterWAV {
    ResourceImporter
}

