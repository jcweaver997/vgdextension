module vgdextension

@[noinit]
pub struct VisualShaderNodeFaceForward {
    VisualShaderNodeVectorBase
}

