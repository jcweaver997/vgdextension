module vgdextension

pub type VSlider = voidptr

