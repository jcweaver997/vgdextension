module vgdextension

pub struct Popup {
    Window
}

