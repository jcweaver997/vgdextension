module vgdextension

pub struct VisualShaderNodeDistanceFade {
    VisualShaderNode
}

