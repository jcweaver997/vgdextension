module vgdextension

pub struct ScriptLanguageExtensionProfilingInfo {
    pub mut:
    signature StringName
    call_count u64
    total_time u64
    self_time u64
}

