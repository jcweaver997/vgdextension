module vgdextension

pub type MovieWriterMJPEG = voidptr

