module vgdextension

pub struct EditorExportPlatformAndroid {
    EditorExportPlatform
}

