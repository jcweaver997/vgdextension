module vgdextension

@[noinit]
pub struct AudioBusLayout {
    Resource
}

