module vgdextension

@[noinit]
pub struct HFlowContainer {
    FlowContainer
}

