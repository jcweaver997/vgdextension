module vgdextension

pub type VBoxContainer = voidptr

