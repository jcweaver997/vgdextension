module vgdextension

pub struct QuadMesh {
    PlaneMesh
}

