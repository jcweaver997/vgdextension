module vgdextension

@[noinit]
pub struct Resource {
    RefCounted
}

pub interface IResourceSetupLocalToScene {
    mut:
    virt_setup_local_to_scene()
}

pub fn (mut r Resource) usetup_local_to_scene() {
    classname := StringName.new("Resource")
    fnname := StringName.new("_setup_local_to_scene")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 0)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (mut r Resource) set_path(path String) {
    classname := StringName.new("Resource")
    fnname := StringName.new("set_path")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 83702148)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&path)}
    gdf.object_method_bind_ptrcall(mb, r.ptr, voidptr(&args[0]), unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (mut r Resource) take_over_path(path String) {
    classname := StringName.new("Resource")
    fnname := StringName.new("take_over_path")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 83702148)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&path)}
    gdf.object_method_bind_ptrcall(mb, r.ptr, voidptr(&args[0]), unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (r &Resource) get_path() String {
    mut object_out := String{}
    classname := StringName.new("Resource")
    fnname := StringName.new("get_path")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 201670096)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, voidptr(&object_out))
    classname.deinit()
    fnname.deinit()
   return object_out
}
pub fn (mut r Resource) set_name(name String) {
    classname := StringName.new("Resource")
    fnname := StringName.new("set_name")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 83702148)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&name)}
    gdf.object_method_bind_ptrcall(mb, r.ptr, voidptr(&args[0]), unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (r &Resource) get_name() String {
    mut object_out := String{}
    classname := StringName.new("Resource")
    fnname := StringName.new("get_name")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 201670096)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, voidptr(&object_out))
    classname.deinit()
    fnname.deinit()
   return object_out
}
pub fn (r &Resource) get_rid() RID {
    mut object_out := RID{}
    classname := StringName.new("Resource")
    fnname := StringName.new("get_rid")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2944877500)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, voidptr(&object_out))
    classname.deinit()
    fnname.deinit()
   return object_out
}
pub fn (mut r Resource) set_local_to_scene(enable bool) {
    classname := StringName.new("Resource")
    fnname := StringName.new("set_local_to_scene")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&enable)}
    gdf.object_method_bind_ptrcall(mb, r.ptr, voidptr(&args[0]), unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (r &Resource) is_local_to_scene() bool {
    mut object_out := false
    classname := StringName.new("Resource")
    fnname := StringName.new("is_local_to_scene")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, voidptr(&object_out))
    classname.deinit()
    fnname.deinit()
   return object_out
}
pub fn (r &Resource) get_local_scene() Node {
    mut object_out := Node{}
    classname := StringName.new("Resource")
    fnname := StringName.new("get_local_scene")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3160264692)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, voidptr(&object_out))
    classname.deinit()
    fnname.deinit()
   return object_out
}
pub fn (mut r Resource) setup_local_to_scene() {
    classname := StringName.new("Resource")
    fnname := StringName.new("setup_local_to_scene")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (mut r Resource) emit_changed() {
    classname := StringName.new("Resource")
    fnname := StringName.new("emit_changed")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
    gdf.object_method_bind_ptrcall(mb, r.ptr, unsafe{nil}, unsafe{nil})
    classname.deinit()
    fnname.deinit()
}
pub fn (r &Resource) duplicate(subresources bool) Resource {
    mut object_out := Resource{}
    classname := StringName.new("Resource")
    fnname := StringName.new("duplicate")
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 482882304)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&subresources)}
    gdf.object_method_bind_ptrcall(mb, r.ptr, voidptr(&args[0]), voidptr(&object_out))
    classname.deinit()
    fnname.deinit()
   return object_out
}
