module vgdextension

pub struct Texture {
    Resource
}

