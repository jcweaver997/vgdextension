module vgdextension

pub struct AnimationNodeTimeScale {
    AnimationNode
}

