module vgdextension

pub type VisualShaderNodeParticleOutput = voidptr

