module vgdextension

pub struct VScrollBar {
    ScrollBar
}

