module vgdextension

@[noinit]
pub struct VisualShaderNodeVectorRefract {
    VisualShaderNodeVectorBase
}

