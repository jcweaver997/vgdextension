module vgdextension

@[noinit]
pub struct CSGCombiner3D {
    CSGShape3D
}

