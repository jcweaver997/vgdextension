module vgdextension

pub struct LightmapperRD {
    Lightmapper
}

