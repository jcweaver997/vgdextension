module vgdextension

pub struct VisualShaderNodeConstant {
    VisualShaderNode
}

