module vgdextension

pub struct SkeletonProfileHumanoid {
    SkeletonProfile
}

