module vgdextension

@[noinit]
pub struct PanelContainer {
    Container
}

