module vgdextension

@[noinit]
pub struct LightmapperRD {
    Lightmapper
}

