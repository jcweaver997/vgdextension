module vgdextension

pub struct AnimationNodeBlend3 {
    AnimationNodeSync
}

