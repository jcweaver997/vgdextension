module vgdextension

pub struct CompressedCubemap {
    CompressedTextureLayered
}

