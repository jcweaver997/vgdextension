module vgdextension

pub type Panel = voidptr

