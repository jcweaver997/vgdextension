module vgdextension

pub struct CheckBox {
    Button
}

