module vgdextension

pub struct TextServerAdvanced {
    TextServerExtension
}

