module vgdextension

@[noinit]
pub struct AnimationNodeAdd3 {
    AnimationNodeSync
}

