module vgdextension

pub struct VisualShaderNodeSDFRaymarch {
    VisualShaderNode
}

