module vgdextension

pub type EditorSceneFormatImporterFBX = voidptr

