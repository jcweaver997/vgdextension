module vgdextension

@[noinit]
pub struct AnimationNodeAdd2 {
    AnimationNodeSync
}

