module vgdextension

pub struct GLTFDocumentExtensionTextureWebP {
    GLTFDocumentExtension
}

