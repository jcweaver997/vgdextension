module vgdextension

pub type AudioEffectLowPassFilter = voidptr

