module vgdextension

@[noinit]
pub struct TextureCubemapArrayRD {
    TextureLayeredRD
}

