module vgdextension

pub struct ORMMaterial3D {
    BaseMaterial3D
}

