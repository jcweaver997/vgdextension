module vgdextension

pub type VisualShaderNodeTexture3DParameter = voidptr

