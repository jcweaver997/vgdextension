module vgdextension

pub type EditorExportPlatformWindows = voidptr

