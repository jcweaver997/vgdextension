module vgdextension

@[noinit]
pub struct ResourceImporterBitMap {
    ResourceImporter
}

