module vgdextension

@[noinit]
pub struct AudioEffectEQ10 {
    AudioEffectEQ
}

