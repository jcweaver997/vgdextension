module vgdextension

pub struct VisualShaderNodeTexture3DParameter {
    VisualShaderNodeTextureParameter
}

