module vgdextension

pub type AnimationNodeAdd2 = voidptr

