module vgdextension

@[noinit]
pub struct AudioEffectEQ21 {
    AudioEffectEQ
}

