module vgdextension

@[noinit]
pub struct PlaceholderTexture2DArray {
    PlaceholderTextureLayered
}

