module vgdextension

pub type VFlowContainer = voidptr

