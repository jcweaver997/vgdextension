module vgdextension

pub type EditorExportPlatformAndroid = voidptr

