module vgdextension

@[noinit]
pub struct IntervalTweener {
    Tweener
}

