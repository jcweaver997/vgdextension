module vgdextension

pub struct OfflineMultiplayerPeer {
    MultiplayerPeer
}

