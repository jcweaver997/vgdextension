module vgdextension

pub struct VisualShaderNodeVaryingSetter {
    VisualShaderNodeVarying
}

