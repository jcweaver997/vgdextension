module vgdextension

pub struct GLTFDocumentExtensionPhysics {
    GLTFDocumentExtension
}

