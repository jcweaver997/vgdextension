module vgdextension

pub struct JavaScriptObject {
    RefCounted
}

