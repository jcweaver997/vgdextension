module vgdextension

@[noinit]
pub struct ShaderGlobalsOverride {
    Node
}

