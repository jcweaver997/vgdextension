module vgdextension

pub struct VisualShaderNodeVaryingGetter {
    VisualShaderNodeVarying
}

