module vgdextension

pub struct VSplitContainer {
    SplitContainer
}

