module vgdextension

@[noinit]
pub struct AudioEffectHighPassFilter {
    AudioEffectFilter
}

