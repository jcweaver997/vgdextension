module vgdextension

pub struct VisualShaderNodeParticleRingEmitter {
    VisualShaderNodeParticleEmitter
}

