module vgdextension

pub type JavaScriptObject = voidptr

