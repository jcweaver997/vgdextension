module vgdextension

@[noinit]
pub struct ResourceImporterTexture {
    ResourceImporter
}

