module vgdextension

pub struct EditorSceneFormatImporterGLTF {
    EditorSceneFormatImporter
}

