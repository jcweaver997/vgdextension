module vgdextension

@[noinit]
pub struct AnimationNodeBlend2 {
    AnimationNodeSync
}

