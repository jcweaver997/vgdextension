module vgdextension

pub type PhysicsDirectBodyState2D = voidptr

pub fn (r &PhysicsDirectBodyState2D) get_total_gravity() Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_total_gravity")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_total_linear_damp() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_total_linear_damp")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_total_angular_damp() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_total_angular_damp")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_center_of_mass() Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_center_of_mass")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_center_of_mass_local() Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_center_of_mass_local")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_inverse_mass() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_inverse_mass")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_inverse_inertia() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_inverse_inertia")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) set_linear_velocity(velocity Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_linear_velocity")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PhysicsDirectBodyState2D) get_linear_velocity() Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_linear_velocity")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) set_angular_velocity(velocity f32) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_angular_velocity")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PhysicsDirectBodyState2D) get_angular_velocity() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_angular_velocity")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) set_transform(transform Transform2D) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_transform")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2761652528)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PhysicsDirectBodyState2D) get_transform() Transform2D {
    mut object_out := Transform2D{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_transform")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3814499831)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_velocity_at_local_position(local_position Vector2) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_velocity_at_local_position")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2656412154)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&local_position)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) apply_central_impulse(impulse Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("apply_central_impulse")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) apply_torque_impulse(impulse f32) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("apply_torque_impulse")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) apply_impulse(impulse Vector2, position Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("apply_impulse")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 496058220)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) apply_central_force(force Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("apply_central_force")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3862383994)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) apply_force(force Vector2, position Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("apply_force")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 496058220)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) apply_torque(torque f32) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("apply_torque")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) add_constant_central_force(force Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("add_constant_central_force")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3862383994)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) add_constant_force(force Vector2, position Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("add_constant_force")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 496058220)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) add_constant_torque(torque f32) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("add_constant_torque")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) set_constant_force(force Vector2) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_constant_force")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 743155724)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PhysicsDirectBodyState2D) get_constant_force() Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_constant_force")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3341600327)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) set_constant_torque(torque f32) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_constant_torque")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PhysicsDirectBodyState2D) get_constant_torque() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_constant_torque")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) set_sleep_state(enabled bool) {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_sleep_state")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2586408642)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PhysicsDirectBodyState2D) is_sleeping() bool {
    mut object_out := false
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("is_sleeping")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 36873697)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_count() i32 {
    mut object_out := i32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_count")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3905245786)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_local_position(contact_idx i32) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_local_position")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2299179447)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_local_normal(contact_idx i32) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_local_normal")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2299179447)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_local_shape(contact_idx i32) i32 {
    mut object_out := i32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_local_shape")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_local_velocity_at_position(contact_idx i32) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_local_velocity_at_position")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2299179447)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_collider(contact_idx i32) RID {
    mut object_out := RID{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_collider")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 495598643)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_collider_position(contact_idx i32) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_collider_position")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2299179447)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_collider_id(contact_idx i32) i32 {
    mut object_out := i32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_collider_id")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_collider_object(contact_idx i32) Object {
    mut object_out := unsafe{nil}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_collider_object")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3332903315)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_collider_shape(contact_idx i32) i32 {
    mut object_out := i32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_collider_shape")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 923996154)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_collider_velocity_at_position(contact_idx i32) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_collider_velocity_at_position")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2299179447)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_contact_impulse(contact_idx i32) Vector2 {
    mut object_out := Vector2{}
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_contact_impulse")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2299179447)
    mut args := unsafe { [1]voidptr{} }
    args[0] = unsafe{voidptr(&contact_idx)}
    gdf.object_method_bind_ptrcall(mb, voidptr(r), voidptr(&args[0]), voidptr(&object_out))
   return object_out
}
pub fn (r &PhysicsDirectBodyState2D) get_step() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_step")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
pub fn (mut r PhysicsDirectBodyState2D) integrate_forces() {
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("integrate_forces")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 3218959716)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (mut r PhysicsDirectBodyState2D) get_space_state() PhysicsDirectSpaceState2D {
    mut object_out := PhysicsDirectSpaceState2D(unsafe{nil})
    classname := StringName.new("PhysicsDirectBodyState2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_space_state")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 2506717822)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
