module vgdextension

@[noinit]
pub struct VisualShaderNodeOutput {
    VisualShaderNode
}

