module vgdextension

@[noinit]
pub struct VisualShaderNodeConstant {
    VisualShaderNode
}

