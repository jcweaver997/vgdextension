module vgdextension

pub enum Orientation as i64 {
    vertical = 1
    horizontal = 0
}
