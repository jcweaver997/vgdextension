module vgdextension

pub type PointMesh = voidptr

