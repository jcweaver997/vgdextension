module vgdextension

pub type PlaceholderTexture2DArray = voidptr

