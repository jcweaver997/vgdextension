module vgdextension

@[noinit]
pub struct PopupPanel {
    Popup
}

