module vgdextension

@[noinit]
pub struct VisualShaderNodeRotationByAxis {
    VisualShaderNode
}

