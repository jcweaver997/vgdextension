module vgdextension

pub enum MouseButtonMask as i64 {
    mouse_button_mask_left = 1
    mouse_button_mask_right = 2
    mouse_button_mask_middle = 4
    mouse_button_mask_mb_xbutton1 = 128
    mouse_button_mask_mb_xbutton2 = 256
}
