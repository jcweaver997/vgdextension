module vgdextension

@[noinit]
pub struct GDScriptEditorTranslationParserPlugin {
    EditorTranslationParserPlugin
}

