module vgdextension

pub struct AudioFrame {
    pub mut:
    left f32
    right f32
}

