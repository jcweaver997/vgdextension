module vgdextension

@[noinit]
pub struct VisualShaderNodeVaryingSetter {
    VisualShaderNodeVarying
}

