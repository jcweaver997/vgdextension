module vgdextension

@[noinit]
pub struct GLTFDocumentExtensionTextureWebP {
    GLTFDocumentExtension
}

