module vgdextension

@[noinit]
pub struct VisualShaderNodeParticleSphereEmitter {
    VisualShaderNodeParticleEmitter
}

