module vgdextension

pub struct EditorExportPlatformMacOS {
    EditorExportPlatform
}

