module vgdextension

pub type GLTFDocumentExtensionTextureWebP = voidptr

