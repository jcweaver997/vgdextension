module vgdextension

pub enum Orientation {
    vertical = 1
    horizontal = 0
}
