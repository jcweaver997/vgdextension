module vgdextension

pub struct GodotPhysicsServer3D {
    PhysicsServer3D
}

