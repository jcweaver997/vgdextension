module vgdextension

pub struct VideoStreamTheora {
    VideoStream
}

