module vgdextension

pub enum JoyButton {
    joy_button_invalid = -1
    joy_button_a = 0
    joy_button_b = 1
    joy_button_x = 2
    joy_button_y = 3
    joy_button_back = 4
    joy_button_guide = 5
    joy_button_start = 6
    joy_button_left_stick = 7
    joy_button_right_stick = 8
    joy_button_left_shoulder = 9
    joy_button_right_shoulder = 10
    joy_button_dpad_up = 11
    joy_button_dpad_down = 12
    joy_button_dpad_left = 13
    joy_button_dpad_right = 14
    joy_button_misc1 = 15
    joy_button_paddle1 = 16
    joy_button_paddle2 = 17
    joy_button_paddle3 = 18
    joy_button_paddle4 = 19
    joy_button_touchpad = 20
    joy_button_sdl_max = 21
    joy_button_max = 128
}
