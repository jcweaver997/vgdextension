module vgdextension

@[noinit]
pub struct AudioEffectNotchFilter {
    AudioEffectFilter
}

