module vgdextension

@[noinit]
pub struct EditorExportPlatformPC {
    EditorExportPlatform
}

