module vgdextension

pub type VisualShaderNodeVectorDistance = voidptr

