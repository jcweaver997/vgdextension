module vgdextension

pub type Node3DGizmo = voidptr

