module vgdextension

pub struct PlaceholderCubemap {
    PlaceholderTextureLayered
}

