module vgdextension

pub type VisualShaderNodeProximityFade = voidptr

