module vgdextension

pub struct EditorSceneFormatImporterFBX {
    EditorSceneFormatImporter
}

