module vgdextension

@[noinit]
pub struct VisualShaderNodeScreenUVToSDF {
    VisualShaderNode
}

