module vgdextension

pub enum VerticalAlignment as i64 {
    vertical_alignment_top = 0
    vertical_alignment_center = 1
    vertical_alignment_bottom = 2
    vertical_alignment_fill = 3
}
