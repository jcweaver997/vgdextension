module vgdextension

@[noinit]
pub struct ResourceImporterCSVTranslation {
    ResourceImporter
}

