module vgdextension

pub type GDScriptEditorTranslationParserPlugin = voidptr

