module vgdextension

pub type CompressedCubemapArray = voidptr

