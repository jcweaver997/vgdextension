module vgdextension

@[noinit]
pub struct AudioEffectBandPassFilter {
    AudioEffectFilter
}

