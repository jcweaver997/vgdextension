module vgdextension

pub type IPUnix = voidptr

