module vgdextension

pub struct VisualShaderNodeVectorDecompose {
    VisualShaderNodeVectorBase
}

