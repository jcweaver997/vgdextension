module vgdextension

pub type VisualShaderNodeVectorCompose = voidptr

