module vgdextension

pub struct OggPacketSequencePlayback {
    RefCounted
}

