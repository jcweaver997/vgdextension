module vgdextension

@[noinit]
pub struct VisualShaderNodeRemap {
    VisualShaderNode
}

