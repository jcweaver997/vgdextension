module vgdextension

@[noinit]
pub struct VisualShaderNodeDistanceFade {
    VisualShaderNode
}

