module vgdextension

@[noinit]
pub struct CompressedCubemapArray {
    CompressedTextureLayered
}

