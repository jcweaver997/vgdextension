module vgdextension

pub struct VisualShaderNodeSDFToScreenUV {
    VisualShaderNode
}

