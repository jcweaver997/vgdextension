module vgdextension

pub type AudioEffectBandPassFilter = voidptr

