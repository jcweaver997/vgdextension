module vgdextension

pub struct HScrollBar {
    ScrollBar
}

