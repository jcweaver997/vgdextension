module vgdextension

pub type HSeparator = voidptr

