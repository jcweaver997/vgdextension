module vgdextension

pub type VisualShaderNodeParticleRingEmitter = voidptr

