module vgdextension

pub type Popup = voidptr

