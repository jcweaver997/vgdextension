module vgdextension

pub struct VisualShaderNodeParticleSphereEmitter {
    VisualShaderNodeParticleEmitter
}

