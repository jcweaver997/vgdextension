module vgdextension

@[noinit]
pub struct VisualShaderNodeParticleBoxEmitter {
    VisualShaderNodeParticleEmitter
}

