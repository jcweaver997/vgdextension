module vgdextension

@[noinit]
pub struct VisualShaderNodeCubemapParameter {
    VisualShaderNodeTextureParameter
}

