module vgdextension

pub type VisualShaderNodeDistanceFade = voidptr

