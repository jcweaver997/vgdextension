module vgdextension

@[noinit]
pub struct VisualShaderNodeTexture2DParameter {
    VisualShaderNodeTextureParameter
}

