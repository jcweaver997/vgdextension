module vgdextension

pub type VisualShaderNodeTextureSDF = voidptr

