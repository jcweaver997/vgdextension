module vgdextension

@[noinit]
pub struct ResourceImporterBMFont {
    ResourceImporter
}

