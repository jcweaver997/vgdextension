module vgdextension

@[noinit]
pub struct VisualShaderNodeTransformCompose {
    VisualShaderNode
}

