module vgdextension

@[noinit]
pub struct Node3DGizmo {
    RefCounted
}

