module vgdextension

pub struct PointMesh {
    PrimitiveMesh
}

