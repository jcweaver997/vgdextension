module vgdextension

pub type ShaderGlobalsOverride = voidptr

