module vgdextension

@[noinit]
pub struct MarginContainer {
    Container
}

