module vgdextension

pub struct VisualShaderNodeLinearSceneDepth {
    VisualShaderNode
}

