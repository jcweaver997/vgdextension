module vgdextension

@[noinit]
pub struct CompressedTexture2DArray {
    CompressedTextureLayered
}

