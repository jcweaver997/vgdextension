module vgdextension

@[noinit]
pub struct EditorSceneFormatImporterBlend {
    EditorSceneFormatImporter
}

