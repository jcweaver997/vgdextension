module vgdextension

pub type VisualShaderNodeConstant = voidptr

