module vgdextension

@[noinit]
pub struct GodotPhysicsServer3D {
    PhysicsServer3D
}

