module vgdextension

pub struct PlaceholderTexture2DArray {
    PlaceholderTextureLayered
}

