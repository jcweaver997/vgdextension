module vgdextension

@[noinit]
pub struct TextServerDummy {
    TextServerExtension
}

