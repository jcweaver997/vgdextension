module vgdextension

pub type AudioEffectBandLimitFilter = voidptr

