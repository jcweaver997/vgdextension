module vgdextension

pub struct Node3DGizmo {
    RefCounted
}

