module vgdextension

@[noinit]
pub struct StandardMaterial3D {
    BaseMaterial3D
}

