module vgdextension

pub type AudioEffectEQ6 = voidptr

