module vgdextension

pub struct HSlider {
    Slider
}

