module vgdextension

@[noinit]
pub struct Texture2DArrayRD {
    TextureLayeredRD
}

