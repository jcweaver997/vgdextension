module vgdextension

pub type CompressedCubemap = voidptr

