module vgdextension

pub enum MouseButton {
    mouse_button_none = 0
    mouse_button_left = 1
    mouse_button_right = 2
    mouse_button_middle = 3
    mouse_button_wheel_up = 4
    mouse_button_wheel_down = 5
    mouse_button_wheel_left = 6
    mouse_button_wheel_right = 7
    mouse_button_xbutton1 = 8
    mouse_button_xbutton2 = 9
}
