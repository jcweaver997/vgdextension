module vgdextension

pub type MarginContainer = voidptr

