module vgdextension

pub type VisualShaderNodeVaryingGetter = voidptr

