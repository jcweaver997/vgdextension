module vgdextension

pub struct VBoxContainer {
    BoxContainer
}

