module vgdextension

@[noinit]
pub struct IPUnix {
    IP
}

