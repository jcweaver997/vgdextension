module vgdextension

@[noinit]
pub struct VisualShaderNodeLinearSceneDepth {
    VisualShaderNode
}

