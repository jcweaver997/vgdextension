module vgdextension

pub struct StyleBoxEmpty {
    StyleBox
}

