module vgdextension

pub type VisualShaderNodeTexture2DParameter = voidptr

