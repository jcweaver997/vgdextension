module vgdextension

pub type VisualShaderNodeFaceForward = voidptr

