module vgdextension

pub type VideoStreamTheora = voidptr

