module vgdextension

@[noinit]
pub struct VSlider {
    Slider
}

