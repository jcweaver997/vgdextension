module vgdextension

pub struct AnimationRootNode {
    AnimationNode
}

