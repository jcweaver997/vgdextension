module vgdextension

pub struct VisualShaderNodeVectorRefract {
    VisualShaderNodeVectorBase
}

