module vgdextension

@[noinit]
pub struct JavaClass {
    RefCounted
}

