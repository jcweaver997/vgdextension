module vgdextension

pub struct PanelContainer {
    Container
}

