module vgdextension

pub struct AnimationNodeBlend2 {
    AnimationNodeSync
}

