module vgdextension

pub struct HSplitContainer {
    SplitContainer
}

