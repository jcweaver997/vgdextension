module vgdextension

pub struct VisualShaderNodeDotProduct {
    VisualShaderNode
}

