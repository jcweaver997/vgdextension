module vgdextension

pub struct Panel {
    Control
}

