module vgdextension

pub type Separator = voidptr

