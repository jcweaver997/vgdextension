module vgdextension

pub type VisualShaderNodeVectorLen = voidptr

