module vgdextension

pub type VisualShaderNodeDeterminant = voidptr

