module vgdextension

pub type VisualShaderNodeCubemapParameter = voidptr

