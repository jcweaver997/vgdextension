module vgdextension

pub struct MovieWriterMJPEG {
    MovieWriter
}

