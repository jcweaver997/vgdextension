module vgdextension

pub type Path3D = voidptr

pub fn (mut r Path3D) set_curve(curve Curve3D) {
    classname := StringName.new("Path3D")
    defer { classname.deinit() }
    fnname := StringName.new("set_curve")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 408955118)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &Path3D) get_curve() Curve3D {
    mut object_out := Curve3D(unsafe{nil})
    classname := StringName.new("Path3D")
    defer { classname.deinit() }
    fnname := StringName.new("get_curve")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 4244715212)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
