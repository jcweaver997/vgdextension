module vgdextension

pub type LightmapProbe = voidptr

