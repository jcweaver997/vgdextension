module vgdextension

@[noinit]
pub struct AudioEffectEQ6 {
    AudioEffectEQ
}

