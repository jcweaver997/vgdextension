module vgdextension

@[noinit]
pub struct VSplitContainer {
    SplitContainer
}

