module vgdextension

pub enum HorizontalAlignment {
    horizontal_alignment_left = 0
    horizontal_alignment_center = 1
    horizontal_alignment_right = 2
    horizontal_alignment_fill = 3
}
