module vgdextension

pub struct AnimationNodeOutput {
    AnimationNode
}

