module vgdextension

pub type PanelContainer = voidptr

