module vgdextension

@[noinit]
pub struct EditorSceneFormatImporterFBX {
    EditorSceneFormatImporter
}

