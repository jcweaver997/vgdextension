module vgdextension

pub struct PhysicsServer2DExtensionRayResult {
    pub mut:
    position Vector2
    normal Vector2
    rid RID
    collider_id ObjectID
    collider &Object
    shape i64
}

