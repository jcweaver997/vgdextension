module vgdextension

pub type MovieWriterPNGWAV = voidptr

