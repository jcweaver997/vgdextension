module vgdextension

@[noinit]
pub struct ResourceImporterImageFont {
    ResourceImporter
}

