module vgdextension

pub struct AudioBusLayout {
    Resource
}

