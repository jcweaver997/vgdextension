module vgdextension

@[noinit]
pub struct JNISingleton {
    Object
}

