module vgdextension

pub struct GLTFDocumentExtensionConvertImporterMesh {
    GLTFDocumentExtension
}

