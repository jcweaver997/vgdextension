module vgdextension

pub enum PropertyHint {
    property_hint_none = 0
    property_hint_range = 1
    property_hint_enum = 2
    property_hint_enum_suggestion = 3
    property_hint_exp_easing = 4
    property_hint_link = 5
    property_hint_flags = 6
    property_hint_layers_2d_render = 7
    property_hint_layers_2d_physics = 8
    property_hint_layers_2d_navigation = 9
    property_hint_layers_3d_render = 10
    property_hint_layers_3d_physics = 11
    property_hint_layers_3d_navigation = 12
    property_hint_layers_avoidance = 37
    property_hint_file = 13
    property_hint_dir = 14
    property_hint_global_file = 15
    property_hint_global_dir = 16
    property_hint_resource_type = 17
    property_hint_multiline_text = 18
    property_hint_expression = 19
    property_hint_placeholder_text = 20
    property_hint_color_no_alpha = 21
    property_hint_object_id = 22
    property_hint_type_string = 23
    property_hint_node_path_to_edited_node = 24
    property_hint_object_too_big = 25
    property_hint_node_path_valid_types = 26
    property_hint_save_file = 27
    property_hint_global_save_file = 28
    property_hint_int_is_objectid = 29
    property_hint_int_is_pointer = 30
    property_hint_array_type = 31
    property_hint_locale_id = 32
    property_hint_localizable_string = 33
    property_hint_node_type = 34
    property_hint_hide_quaternion_edit = 35
    property_hint_password = 36
    property_hint_max = 38
}
