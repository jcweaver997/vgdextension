module vgdextension

pub enum Corner as i64 {
    corner_top_left = 0
    corner_top_right = 1
    corner_bottom_right = 2
    corner_bottom_left = 3
}
