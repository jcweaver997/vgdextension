module vgdextension

pub type AudioEffectEQ21 = voidptr

