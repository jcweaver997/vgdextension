module vgdextension

@[noinit]
pub struct VisualShaderNodeUVPolarCoord {
    VisualShaderNode
}

