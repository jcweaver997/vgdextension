module vgdextension

@[noinit]
pub struct VisualShaderNodeParticleConeVelocity {
    VisualShaderNode
}

