module vgdextension

pub type JNISingleton = voidptr

