module vgdextension

pub struct IPUnix {
    IP
}

