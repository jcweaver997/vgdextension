module vgdextension

@[noinit]
pub struct VisualShaderNodeVectorLen {
    VisualShaderNodeVectorBase
}

