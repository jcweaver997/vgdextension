module vgdextension

pub type VisualShaderNodeTransformCompose = voidptr

