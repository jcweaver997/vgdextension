module vgdextension

pub type AnimationNodeBlend2 = voidptr

