module vgdextension

pub struct StandardMaterial3D {
    BaseMaterial3D
}

