module vgdextension

@[noinit]
pub struct VSeparator {
    Separator
}

