module vgdextension

pub type StandardMaterial3D = voidptr

