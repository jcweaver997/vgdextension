module vgdextension

@[noinit]
pub struct ResourceFormatImporterSaver {
    ResourceFormatSaver
}

