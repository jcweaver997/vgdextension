module vgdextension

pub struct AudioEffectLowPassFilter {
    AudioEffectFilter
}

