module vgdextension

pub struct XRCamera3D {
    Camera3D
}

