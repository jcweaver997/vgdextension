module vgdextension

pub struct ShaderGlobalsOverride {
    Node
}

