module vgdextension

pub type SkeletonProfileHumanoid = voidptr

