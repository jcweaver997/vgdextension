module vgdextension

pub struct VisualShaderNodeParticleOutput {
    VisualShaderNodeOutput
}

