module vgdextension

@[noinit]
pub struct EditorExportPlatformIOS {
    EditorExportPlatform
}

