module vgdextension

@[noinit]
pub struct MovieWriterPNGWAV {
    MovieWriter
}

