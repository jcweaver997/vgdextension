module vgdextension

@[noinit]
pub struct VisualShaderNodeTextureParameterTriplanar {
    VisualShaderNodeTextureParameter
}

