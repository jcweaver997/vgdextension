module vgdextension

pub type AudioBusLayout = voidptr

