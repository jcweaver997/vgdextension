module vgdextension

pub type AudioEffectLowShelfFilter = voidptr

