module vgdextension

@[noinit]
pub struct OggPacketSequencePlayback {
    RefCounted
}

