module vgdextension

@[noinit]
pub struct VisualShaderNodeVaryingGetter {
    VisualShaderNodeVarying
}

