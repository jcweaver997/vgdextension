module vgdextension

pub type VisualShaderNodeVectorDecompose = voidptr

