module vgdextension

@[noinit]
pub struct PlaceholderCubemapArray {
    PlaceholderTextureLayered
}

