module vgdextension

@[noinit]
pub struct CheckBox {
    Button
}

