module vgdextension

pub struct VisualShaderNodeGlobalExpression {
    VisualShaderNodeExpression
}

