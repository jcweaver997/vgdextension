module vgdextension

pub type VisualShaderNodeSDFToScreenUV = voidptr

