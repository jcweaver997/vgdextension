module vgdextension

pub struct Separator {
    Control
}

