module vgdextension

@[noinit]
pub struct MovieWriterMJPEG {
    MovieWriter
}

