module vgdextension

pub enum EulerOrder {
    euler_order_xyz = 0
    euler_order_xzy = 1
    euler_order_yxz = 2
    euler_order_yzx = 3
    euler_order_zxy = 4
    euler_order_zyx = 5
}
