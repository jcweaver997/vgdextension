module vgdextension

pub type AnimationNodeBlend3 = voidptr

