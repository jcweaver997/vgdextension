module vgdextension

pub type AudioEffectHighPassFilter = voidptr

