module vgdextension

pub type VisualShaderNodeParticleSphereEmitter = voidptr

