module vgdextension

pub type GodotPhysicsServer3D = voidptr

