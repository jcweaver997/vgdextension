module vgdextension

pub type VisualShaderNodeUVPolarCoord = voidptr

