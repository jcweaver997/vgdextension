module vgdextension

@[noinit]
pub struct Panel {
    Control
}

