module vgdextension

pub struct VisualShaderNodeVectorDistance {
    VisualShaderNodeVectorBase
}

