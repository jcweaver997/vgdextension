module vgdextension

@[noinit]
pub struct ORMMaterial3D {
    BaseMaterial3D
}

