module vgdextension

@[noinit]
pub struct VisualShaderNodeScreenNormalWorldSpace {
    VisualShaderNode
}

