module vgdextension

pub struct AudioEffectLowShelfFilter {
    AudioEffectFilter
}

