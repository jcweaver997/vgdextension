module vgdextension

pub struct GDScriptEditorTranslationParserPlugin {
    EditorTranslationParserPlugin
}

