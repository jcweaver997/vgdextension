module vgdextension

@[noinit]
pub struct ResourceImporterTextureAtlas {
    ResourceImporter
}

