module vgdextension

@[noinit]
pub struct VisualShaderNodeFresnel {
    VisualShaderNode
}

