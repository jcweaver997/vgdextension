module vgdextension

pub type OggPacketSequencePlayback = voidptr

