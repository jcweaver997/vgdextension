module vgdextension

pub struct VisualShaderNodeParticleBoxEmitter {
    VisualShaderNodeParticleEmitter
}

