module vgdextension

@[noinit]
pub struct CompressedCubemap {
    CompressedTextureLayered
}

