module vgdextension

pub struct MarginContainer {
    Container
}

