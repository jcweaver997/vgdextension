module vgdextension

pub type VisualShaderNodeSDFRaymarch = voidptr

