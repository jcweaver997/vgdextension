module vgdextension

pub type VisualShaderNodeParticleConeVelocity = voidptr

