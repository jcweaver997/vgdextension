module vgdextension

pub struct JNISingleton {
    Object
}

