module vgdextension

pub struct VisualShaderNodeTextureSDF {
    VisualShaderNode
}

