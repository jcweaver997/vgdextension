module vgdextension

pub struct AudioEffectBandLimitFilter {
    AudioEffectFilter
}

