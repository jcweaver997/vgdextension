module vgdextension

@[noinit]
pub struct AnimationNodeTimeSeek {
    AnimationNode
}

