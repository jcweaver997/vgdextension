module vgdextension

pub type AnimationRootNode = voidptr

