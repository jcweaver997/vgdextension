module vgdextension

pub struct HBoxContainer {
    BoxContainer
}

