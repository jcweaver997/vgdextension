module vgdextension

pub type HSlider = voidptr

