module vgdextension

pub struct PopupPanel {
    Popup
}

