module vgdextension

@[noinit]
pub struct VFlowContainer {
    FlowContainer
}

