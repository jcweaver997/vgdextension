module vgdextension

pub type EditorSceneFormatImporterBlend = voidptr

