module vgdextension

@[noinit]
pub struct VisualShaderNodeVectorDistance {
    VisualShaderNodeVectorBase
}

