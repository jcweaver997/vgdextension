module vgdextension

pub struct VisualShaderNodeOutput {
    VisualShaderNode
}

