module vgdextension

@[noinit]
pub struct VisualShaderNodeSDFRaymarch {
    VisualShaderNode
}

