module vgdextension

@[noinit]
pub struct VisualShaderNodeTransformDecompose {
    VisualShaderNode
}

