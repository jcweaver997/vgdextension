module vgdextension

pub struct VSlider {
    Slider
}

