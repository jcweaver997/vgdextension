module vgdextension

pub type VisualShaderNodeTextureSDFNormal = voidptr

