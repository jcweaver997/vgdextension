module vgdextension

pub type EditorExportPlatformLinuxBSD = voidptr

