module vgdextension

pub enum ClockDirection as i64 {
    clockwise = 0
    counterclockwise = 1
}
