module vgdextension

@[noinit]
pub struct VideoStreamTheora {
    VideoStream
}

