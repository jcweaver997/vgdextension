module vgdextension

pub type PlaceholderCubemapArray = voidptr

