module vgdextension

@[noinit]
pub struct AudioEffectLowShelfFilter {
    AudioEffectFilter
}

