module vgdextension

pub type StyleBoxEmpty = voidptr

