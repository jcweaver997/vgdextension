module vgdextension

pub struct VisualShaderNodeRemap {
    VisualShaderNode
}

