module vgdextension

pub type PinJoint2D = voidptr

pub fn (mut r PinJoint2D) set_softness(softness f32) {
    classname := StringName.new("PinJoint2D")
    defer { classname.deinit() }
    fnname := StringName.new("set_softness")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &PinJoint2D) get_softness() f32 {
    mut object_out := f32(0)
    classname := StringName.new("PinJoint2D")
    defer { classname.deinit() }
    fnname := StringName.new("get_softness")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
