module vgdextension

pub struct VisualShaderNodeTexture2DParameter {
    VisualShaderNodeTextureParameter
}

