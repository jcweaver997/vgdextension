module vgdextension

pub enum JoyAxis {
    joy_axis_invalid = -1
    joy_axis_left_x = 0
    joy_axis_left_y = 1
    joy_axis_right_x = 2
    joy_axis_right_y = 3
    joy_axis_trigger_left = 4
    joy_axis_trigger_right = 5
    joy_axis_sdl_max = 6
    joy_axis_max = 10
}
