module vgdextension

pub struct HSeparator {
    Separator
}

