module vgdextension

@[noinit]
pub struct AudioEffectBandLimitFilter {
    AudioEffectFilter
}

