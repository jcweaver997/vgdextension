module vgdextension

pub type EditorExportPlatformPC = voidptr

