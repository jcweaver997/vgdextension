module vgdextension

pub struct Lightmapper {
    RefCounted
}

