module vgdextension

pub type AudioEffectHighShelfFilter = voidptr

