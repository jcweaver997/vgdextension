module vgdextension

pub struct AnimationNodeTimeSeek {
    AnimationNode
}

