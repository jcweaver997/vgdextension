module vgdextension

pub type XRCamera3D = voidptr

