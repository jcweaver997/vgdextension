module vgdextension

pub struct AudioEffectHighPassFilter {
    AudioEffectFilter
}

