module vgdextension

@[noinit]
pub struct AudioEffectHighShelfFilter {
    AudioEffectFilter
}

