module vgdextension

pub enum MethodFlags {
    method_flag_normal = 1
    method_flag_editor = 2
    method_flag_const = 4
    method_flag_virtual = 8
    method_flag_vararg = 16
    method_flag_static = 32
    method_flag_object_core = 64
}
