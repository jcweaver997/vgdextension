module vgdextension

@[noinit]
pub struct JavaScriptObject {
    RefCounted
}

