module vgdextension

pub type PlaceholderCubemap = voidptr

