module vgdextension

pub struct TextServerDummy {
    TextServerExtension
}

