module vgdextension

pub type VisualShaderNodeRandomRange = voidptr

