module vgdextension

pub struct EditorExportPlatform {
    RefCounted
}

