module vgdextension

@[noinit]
pub struct PointMesh {
    PrimitiveMesh
}

