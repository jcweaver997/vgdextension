module vgdextension

pub struct PlaceholderMaterial {
    Material
}

