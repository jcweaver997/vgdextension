module vgdextension

pub type VisualShaderNodeIf = voidptr

