module vgdextension

pub type CheckButton = voidptr

