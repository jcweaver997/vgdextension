module vgdextension

pub type TextServerAdvanced = voidptr

