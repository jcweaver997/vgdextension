module vgdextension

pub type AnimationNodeSub2 = voidptr

