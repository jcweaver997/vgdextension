module vgdextension

@[noinit]
pub struct XRCamera3D {
    Camera3D
}

