module vgdextension

pub type VisualShaderNodeTexture2DArrayParameter = voidptr

