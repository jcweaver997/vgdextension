module vgdextension

pub enum VariantType as i64 {
    type_nil = 0
    type_bool = 1
    type_int = 2
    type_float = 3
    type_string = 4
    type_vector2 = 5
    type_vector2i = 6
    type_rect2 = 7
    type_rect2i = 8
    type_vector3 = 9
    type_vector3i = 10
    type_transform2d = 11
    type_vector4 = 12
    type_vector4i = 13
    type_plane = 14
    type_quaternion = 15
    type_aabb = 16
    type_basis = 17
    type_transform3d = 18
    type_projection = 19
    type_color = 20
    type_string_name = 21
    type_node_path = 22
    type_rid = 23
    type_object = 24
    type_callable = 25
    type_signal = 26
    type_dictionary = 27
    type_array = 28
    type_packed_byte_array = 29
    type_packed_int32_array = 30
    type_packed_int64_array = 31
    type_packed_float32_array = 32
    type_packed_float64_array = 33
    type_packed_string_array = 34
    type_packed_vector2_array = 35
    type_packed_vector3_array = 36
    type_packed_color_array = 37
    type_max = 38
}
