module vgdextension

@[noinit]
pub struct Texture {
    Resource
}

