module vgdextension

@[noinit]
pub struct VisualShaderNodeParticleRingEmitter {
    VisualShaderNodeParticleEmitter
}

