module vgdextension

@[noinit]
pub struct ResourceImporterDynamicFont {
    ResourceImporter
}

