module vgdextension

pub type HFlowContainer = voidptr

