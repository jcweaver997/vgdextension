module vgdextension

pub type AnimationNodeOutput = voidptr

