module vgdextension

pub type VisualShaderNodeDotProduct = voidptr

