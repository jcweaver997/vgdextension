module vgdextension

pub struct VisualShaderNodeFresnel {
    VisualShaderNode
}

