module vgdextension

pub type VSeparator = voidptr

