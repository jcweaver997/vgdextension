module vgdextension

pub type AnimationNodeAdd3 = voidptr

