module vgdextension

pub type Lightmapper = voidptr

