module vgdextension

pub struct VisualShaderNodeTextureParameterTriplanar {
    VisualShaderNodeTextureParameter
}

