module vgdextension

@[noinit]
pub struct AudioStreamMicrophone {
    AudioStream
}

