module vgdextension

pub enum Side as i64 {
    side_left = 0
    side_top = 1
    side_right = 2
    side_bottom = 3
}
