module vgdextension

pub type TriangleMesh = voidptr

