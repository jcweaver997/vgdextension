module vgdextension

@[noinit]
pub struct StyleBoxEmpty {
    StyleBox
}

