module vgdextension

pub struct EditorExportPlatformIOS {
    EditorExportPlatform
}

