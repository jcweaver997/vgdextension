module vgdextension

pub struct AudioStreamMicrophone {
    AudioStream
}

