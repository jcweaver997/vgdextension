module vgdextension

pub struct TriangleMesh {
    RefCounted
}

