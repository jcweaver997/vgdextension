module vgdextension

pub struct VisualShaderNodeProximityFade {
    VisualShaderNode
}

