module vgdextension

pub type HSplitContainer = voidptr

