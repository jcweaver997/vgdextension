module vgdextension

@[noinit]
pub struct AnimationNodeTimeScale {
    AnimationNode
}

