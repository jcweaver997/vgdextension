module vgdextension

pub struct PhysicsServer3DExtensionShapeResult {
    pub mut:
    rid RID
    collider_id ObjectID
    collider &Object
    shape int
}

