module vgdextension

@[noinit]
pub struct GLTFDocumentExtensionConvertImporterMesh {
    GLTFDocumentExtension
}

