module vgdextension

pub struct VisualShaderNodeTexture2DArrayParameter {
    VisualShaderNodeTextureParameter
}

