module vgdextension

pub struct HFlowContainer {
    FlowContainer
}

