module vgdextension

@[noinit]
pub struct ResourceImporterLayeredTexture {
    ResourceImporter
}

