module vgdextension

pub struct AnimationNodeAdd2 {
    AnimationNodeSync
}

