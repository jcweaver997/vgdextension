module vgdextension

@[noinit]
pub struct EditorExportPlatformMacOS {
    EditorExportPlatform
}

