module vgdextension

pub type VisualShaderNodeRemap = voidptr

