module vgdextension

pub struct VisualShaderNodeOuterProduct {
    VisualShaderNode
}

