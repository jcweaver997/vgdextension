module vgdextension

pub struct JavaClass {
    RefCounted
}

