module vgdextension

pub type TextServerDummy = voidptr

