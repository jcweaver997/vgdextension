module vgdextension

pub struct VisualShaderNodeTransformCompose {
    VisualShaderNode
}

