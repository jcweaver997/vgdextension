module vgdextension

@[noinit]
pub struct ScriptLanguage {
    Object
}

