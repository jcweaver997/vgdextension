module vgdextension

pub type VisualShaderNodeOutput = voidptr

