module vgdextension

@[noinit]
pub struct Lightmapper {
    RefCounted
}

