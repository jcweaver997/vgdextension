module vgdextension

@[noinit]
pub struct VisualShaderNodeTexture2DArrayParameter {
    VisualShaderNodeTextureParameter
}

