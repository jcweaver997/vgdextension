module vgdextension

pub type ResourceFormatImporterSaver = voidptr

