module vgdextension

@[noinit]
pub struct VBoxContainer {
    BoxContainer
}

