module vgdextension

pub struct PlaceholderCubemapArray {
    PlaceholderTextureLayered
}

