module vgdextension

pub struct ObjectID {
    pub mut:
    id u64
}

