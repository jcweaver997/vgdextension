module vgdextension

@[noinit]
pub struct EditorExportPlatformWindows {
    EditorExportPlatformPC
}

