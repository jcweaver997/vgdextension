module vgdextension

pub type CheckBox = voidptr

