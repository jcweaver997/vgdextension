module vgdextension

pub struct CheckButton {
    Button
}

