module vgdextension

pub struct VisualShaderNodeVectorCompose {
    VisualShaderNodeVectorBase
}

