module vgdextension

@[noinit]
pub struct VisualShaderNodeGlobalExpression {
    VisualShaderNodeExpression
}

