module vgdextension

pub type GPUParticlesCollisionSphere3D = voidptr

pub fn (mut r GPUParticlesCollisionSphere3D) set_radius(radius f32) {
    classname := StringName.new("GPUParticlesCollisionSphere3D")
    defer { classname.deinit() }
    fnname := StringName.new("set_radius")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 373806689)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, unsafe{nil})
}
pub fn (r &GPUParticlesCollisionSphere3D) get_radius() f32 {
    mut object_out := f32(0)
    classname := StringName.new("GPUParticlesCollisionSphere3D")
    defer { classname.deinit() }
    fnname := StringName.new("get_radius")
    defer { fnname.deinit() }
    mb := gdf.classdb_get_method_bind(&classname, &fnname, 1740695150)
    gdf.object_method_bind_ptrcall(mb, voidptr(r), unsafe{nil}, voidptr(&object_out))
   return object_out
}
