module vgdextension

pub type VisualShaderNodeFresnel = voidptr

