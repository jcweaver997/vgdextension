module vgdextension

pub type VSplitContainer = voidptr

