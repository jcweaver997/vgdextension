module vgdextension

pub enum KeyModifierMask {
    key_code_mask = 8388607
    key_modifier_mask = 532676608
    key_mask_cmd_or_ctrl = 16777216
    key_mask_shift = 33554432
    key_mask_alt = 67108864
    key_mask_meta = 134217728
    key_mask_ctrl = 268435456
    key_mask_kpad = 536870912
    key_mask_group_switch = 1073741824
}
