module vgdextension

pub type VScrollBar = voidptr

