module vgdextension

@[noinit]
pub struct TextureCubemapRD {
    TextureLayeredRD
}

