module vgdextension

@[noinit]
pub struct VisualShaderNodeRandomRange {
    VisualShaderNode
}

