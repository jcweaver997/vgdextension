module vgdextension

@[noinit]
pub struct VisualShaderNodeWorldPositionFromDepth {
    VisualShaderNode
}

