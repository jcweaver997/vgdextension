module vgdextension

pub type EditorExportPlatform = voidptr

