module vgdextension

pub type AudioStreamPlaybackOggVorbis = voidptr

