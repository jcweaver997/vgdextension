module vgdextension

@[noinit]
pub struct EditorExportPlatformWeb {
    EditorExportPlatform
}

