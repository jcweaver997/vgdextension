module vgdextension

@[noinit]
pub struct OfflineMultiplayerPeer {
    MultiplayerPeer
}

