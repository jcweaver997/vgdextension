module vgdextension

@[noinit]
pub struct GodotPhysicsServer2D {
    PhysicsServer2D
}

