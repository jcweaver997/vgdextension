module vgdextension

pub type AudioEffectEQ10 = voidptr

