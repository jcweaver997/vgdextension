module vgdextension

pub struct AudioStreamPlaybackOggVorbis {
    AudioStreamPlaybackResampled
}

