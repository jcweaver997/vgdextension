module vgdextension

pub struct EditorExportPlatformWindows {
    EditorExportPlatformPC
}

