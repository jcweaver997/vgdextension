module vgdextension

pub struct AudioEffectEQ21 {
    AudioEffectEQ
}

