module vgdextension

pub struct AnimationNodeAdd3 {
    AnimationNodeSync
}

