module vgdextension

pub struct ResourceFormatImporterSaver {
    ResourceFormatSaver
}

