module vgdextension

pub struct VisualShaderNodeTransformDecompose {
    VisualShaderNode
}

