module vgdextension

pub type GodotPhysicsServer2D = voidptr

