module vgdextension

pub struct AnimationNodeSub2 {
    AnimationNodeSync
}

