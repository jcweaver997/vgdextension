module vgdextension

@[noinit]
pub struct Popup {
    Window
}

