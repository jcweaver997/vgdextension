module vgdextension

@[noinit]
pub struct AnimationRootNode {
    AnimationNode
}

