module vgdextension

pub struct CompressedTexture2DArray {
    CompressedTextureLayered
}

