module vgdextension

@[noinit]
pub struct EditorExportPlatformAndroid {
    EditorExportPlatform
}

