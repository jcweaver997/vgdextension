module vgdextension

@[noinit]
pub struct GLTFDocumentExtensionPhysics {
    GLTFDocumentExtension
}

