module vgdextension

pub struct VisualShaderNodeUVPolarCoord {
    VisualShaderNode
}

