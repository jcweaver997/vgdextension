module vgdextension

@[noinit]
pub struct VisualShaderNodeOuterProduct {
    VisualShaderNode
}

