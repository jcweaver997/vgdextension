module vgdextension

pub struct VisualShaderNodeVectorLen {
    VisualShaderNodeVectorBase
}

