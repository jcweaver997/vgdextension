module vgdextension

@[noinit]
pub struct LightmapProbe {
    Node3D
}

