module vgdextension

pub type Texture = voidptr

