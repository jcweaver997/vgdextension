module vgdextension

pub struct AudioEffectEQ6 {
    AudioEffectEQ
}

