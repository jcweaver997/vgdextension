module vgdextension

pub type PlaceholderMaterial = voidptr

