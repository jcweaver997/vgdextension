module vgdextension

pub enum VerticalAlignment {
    vertical_alignment_top = 0
    vertical_alignment_center = 1
    vertical_alignment_bottom = 2
    vertical_alignment_fill = 3
}
