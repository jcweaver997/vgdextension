module vgdextension

pub struct EditorExportPlatformWeb {
    EditorExportPlatform
}

