module vgdextension

pub struct VSeparator {
    Separator
}

