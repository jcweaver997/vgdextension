module vgdextension

pub struct VisualShaderNodeDeterminant {
    VisualShaderNode
}

