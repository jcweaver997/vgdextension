module vgdextension

@[noinit]
pub struct HSplitContainer {
    SplitContainer
}

