module vgdextension

@[noinit]
pub struct CheckButton {
    Button
}

