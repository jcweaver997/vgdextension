module vgdextension

pub type VisualShaderNodeOuterProduct = voidptr

