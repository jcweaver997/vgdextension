module vgdextension

pub struct ScriptLanguage {
    Object
}

