module vgdextension

@[noinit]
pub struct VisualShaderNodeIf {
    VisualShaderNode
}

