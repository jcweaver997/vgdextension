module vgdextension

pub type PopupPanel = voidptr

