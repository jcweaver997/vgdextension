module vgdextension

pub enum VariantOperator {
    op_equal = 0
    op_not_equal = 1
    op_less = 2
    op_less_equal = 3
    op_greater = 4
    op_greater_equal = 5
    op_add = 6
    op_subtract = 7
    op_multiply = 8
    op_divide = 9
    op_negate = 10
    op_positive = 11
    op_module = 12
    op_power = 13
    op_shift_left = 14
    op_shift_right = 15
    op_bit_and = 16
    op_bit_or = 17
    op_bit_xor = 18
    op_bit_negate = 19
    op_and = 20
    op_or = 21
    op_xor = 22
    op_not = 23
    op_in = 24
    op_max = 25
}
