module vgdextension

@[noinit]
pub struct Tweener {
    RefCounted
}

