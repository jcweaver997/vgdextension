module vgdextension

@[noinit]
pub struct SkeletonProfileHumanoid {
    SkeletonProfile
}

