module vgdextension

pub struct IntervalTweener {
    Tweener
}

