module vgdextension

pub struct GDScript {
    Script
}

