module vgdextension

@[noinit]
pub struct VisualShaderNodeVectorCompose {
    VisualShaderNodeVectorBase
}

