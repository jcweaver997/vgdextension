module vgdextension

pub struct SpotLight3D {
    Light3D
}

