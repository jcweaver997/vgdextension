module vgdextension

@[noinit]
pub struct VisualShaderNodeDotProduct {
    VisualShaderNode
}

