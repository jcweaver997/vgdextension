module vgdextension

pub struct AudioEffectHighShelfFilter {
    AudioEffectFilter
}

