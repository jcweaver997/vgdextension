module vgdextension

pub type GDScript = voidptr

