module vgdextension

pub struct AudioEffectEQ10 {
    AudioEffectEQ
}

