module vgdextension

pub type VisualShaderNodeParticleBoxEmitter = voidptr

