module vgdextension

@[noinit]
pub struct HBoxContainer {
    BoxContainer
}

