module vgdextension

@[noinit]
pub struct ResourceImporterImage {
    ResourceImporter
}

