module vgdextension

pub type GLTFDocumentExtensionConvertImporterMesh = voidptr

