module vgdextension

pub type HScrollBar = voidptr

