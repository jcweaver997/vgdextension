module vgdextension

@[noinit]
pub struct TriangleMesh {
    RefCounted
}

