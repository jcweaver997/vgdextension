module vgdextension

pub struct VisualShaderNodeFaceForward {
    VisualShaderNodeVectorBase
}

