module vgdextension

pub type VisualShaderNodeTextureParameterTriplanar = voidptr

