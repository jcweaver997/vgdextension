module vgdextension

@[noinit]
pub struct PlaceholderMaterial {
    Material
}

