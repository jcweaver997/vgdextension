module vgdextension

pub struct VisualShaderNodeParticleConeVelocity {
    VisualShaderNode
}

