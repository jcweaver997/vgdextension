module vgdextension

pub struct VisualShaderNodeScreenUVToSDF {
    VisualShaderNode
}

