module vgdextension

@[noinit]
pub struct ResourceImporterMP3 {
    ResourceImporter
}

