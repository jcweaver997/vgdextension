module vgdextension

pub type AnimationNodeTimeScale = voidptr

