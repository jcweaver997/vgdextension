module vgdextension

@[noinit]
pub struct VisualShaderNodeDeterminant {
    VisualShaderNode
}

