module vgdextension

pub type VisualShaderNodeTransformDecompose = voidptr

