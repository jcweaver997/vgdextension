module vgdextension

@[noinit]
pub struct HSeparator {
    Separator
}

