module vgdextension

pub struct AudioFrame {
    pub mut:
    left f64
    right f64
}

