module vgdextension

@[noinit]
pub struct QuadMesh {
    PlaneMesh
}

